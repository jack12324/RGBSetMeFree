module FPURequestBufferMemory #(BANK_WIDTH = 8, MEM_BUFFER_DEPTH_BYTES = 512)(wr, clk, rst_n, data_in, write_sel, address, data_out);
endmodule
