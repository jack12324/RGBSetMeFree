module fpu_cache (
    ports
);
    
endmodule