// ***************************************************************************
// Copyright (c) 2017, Intel Corporation
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// * Redistributions of source code must retain the above copyright notice,
// this list of conditions and the following disclaimer.
// * Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
// * Neither the name of Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//
// ***************************************************************************

// ===========================================
// Module to Register SR <--> PR signals in SR
// TODO_START
// Include HSSI ethernet IF
// TODO_END -- Narayanan
// ===========================================

import ccip_if_pkg::*;
module ccip_interface_reg(
  // CCI-P Clocks and Resets
  input           logic             pClk,                    // 400MHz - CC-P clock domain. Primary Clock
  input           logic             pck_cp2af_softReset_T0,  // CCI-P ACTIVE HIGH Soft Reset
  input           logic [1:0]       pck_cp2af_pwrState_T0,   // CCI-P AFU Power State
  input           logic             pck_cp2af_error_T0,      // CCI-P Protocol Error Detected
  // Interface structures
  input           t_if_ccip_Rx      pck_cp2af_sRx_T0,        // CCI-P Rx Port
  input           t_if_ccip_Tx      pck_af2cp_sTx_T0,        // CCI-P Tx Port
  
  output          logic             pck_cp2af_softReset_T1,
  output          logic [1:0]       pck_cp2af_pwrState_T1, 
  output          logic             pck_cp2af_error_T1,    
                                    
  output          t_if_ccip_Rx      pck_cp2af_sRx_T1,      
  output          t_if_ccip_Tx      pck_af2cp_sTx_T1

);
(* preserve *) logic             pck_cp2af_softReset_T0_q;
(* preserve *) logic [1:0]       pck_cp2af_pwrState_T0_q;
(* preserve *) logic             pck_cp2af_error_T0_q;
(* preserve *) t_if_ccip_Rx      pck_cp2af_sRx_T0_q;     
(* preserve *) t_if_ccip_Tx      pck_af2cp_sTx_T0_q;

always@(posedge pClk)
begin
    pck_cp2af_softReset_T0_q   <= pck_cp2af_softReset_T0;
    pck_cp2af_pwrState_T0_q    <= pck_cp2af_pwrState_T0;
    pck_cp2af_error_T0_q       <= pck_cp2af_error_T0;
    pck_cp2af_sRx_T0_q         <= pck_cp2af_sRx_T0;
    pck_af2cp_sTx_T0_q         <= pck_af2cp_sTx_T0;
end

always_comb
begin
    pck_cp2af_softReset_T1      = pck_cp2af_softReset_T0_q;
    pck_cp2af_pwrState_T1       = pck_cp2af_pwrState_T0_q;
    pck_cp2af_error_T1          = pck_cp2af_error_T0_q;
    pck_cp2af_sRx_T1            = pck_cp2af_sRx_T0_q;
    pck_af2cp_sTx_T1            = pck_af2cp_sTx_T0_q;
end

endmodule
