module cpu_cache_ctrl (
    ports
);
    
endmodule