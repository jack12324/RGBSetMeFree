module fpu_cache_ctrl (
    
);
    
endmodule