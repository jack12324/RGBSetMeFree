module fpu_cache_ctrl (
    ports
);
    
endmodule